`define CMD_READ   2'b00
`define CMD_WRITE  2'b01
`define CMD_WREN   2'b10