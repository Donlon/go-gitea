`define JUDGER_INVALID 2'b00
`define JUDGER_VALID   2'b01
`define JUDGER_WIN     2'b10
