`define SIDE_GREEN   1'b0
`define SIDE_RED     1'b1